Alberto //NAME
2       //LVL
3       //XP
15      //GOLD
100     //HP
100     //MaxHP
10      //ATT
10      //DEF
10      //SPE
1       //LUCK
10      //TRINKET ID
11E     //TRINKET EQUIPPED ID
99      //SEP?
00      //CONSUMABLE ID
01      //CONSUMABLE ID
01U2    //CONSUMABLE USED ID USES REMAINING